`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/11/17 17:17:12
// Design Name: 
// Module Name: x4_7seg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/*4λ7�����������ԭ��ÿ��ѡͨ1λ����ʾ��Ӧ���֣�һ��ʱ���ѡͨ��һλ��ʾ��Ӧ���֣�ʱ����ѡ�����ʱ���۹۲쵽���������־��������ġ��������ظ�����
ѡ�����ʱ�伴Ϊ�߶�����ܵķ�Ƶ���⣬Ƶ��̫��(����4λ����ʱ�䳬��20ms)����ܻ������˸����Ƶ��̫�߻��������̫�������޷����壬���һ��ɨ����Ϊ��ms
���ϣ��������̲�����0.02s�������������0.02/4=0.005s����Ƶ����С����Ϊ1/0.005=200Hz
���⣬����һֻ����ܺ���ŵ�ڶ�ֻ����ǰ��Ҫ�ضϵ�һֻ����ܣ��������ֻ���
�˴�����Ƶ��Ϊ400Hz����ʱ���źŵļ�������Ӧȡ(1/400)s / (1/100M)s = 250000����2**18=262144����[17:0]����1�������ж�clk_cnt[19:18]��4��ȡֵ���ɡ�
*/
module x4_7seg(x,clk,a_to_g,an,dp);
    input [15:0] x;         //����4λʮ���������֣��ֱ����ĸ����������ʾ
    input clk;              //clk��ϵͳĬ��ʱ���źţ�Ƶ��Ϊ100MHz
    output reg [6:0]a_to_g; //a_to_g��ʾ�����������ʾ������
    output reg [3:0]an;     //an��ʹ���źţ���ʾ4���������һ��������
    output dp;              //dp��ʾС����
    
    wire [1:0] s;           //��ʱ��������ʾclk_cnt�����λ��4��ֵ�������Ӧan��4��ѡ��
    reg [3:0] digit;        //��ʱ��������ʾ����ʾ��1λ16������
    reg [19:0] clk_cnt=0;   //������������¼clk�仯����
    assign dp=1;
    assign s=clk_cnt[19:18];
    //���¼���always���Ϊ����ִ��
    always@(*)              //ȷ��λ
    case(s)
        2'b00:digit=x[3:0];
        2'b01:digit=x[7:4];
        2'b10:digit=x[11:8];
        2'b11:digit=x[15:12];
        default:digit=x[3:0];
    endcase
    always@(*)              //ȷ��λ
    case(digit)
        4'h0:a_to_g=7'b0000001;
        4'h1:a_to_g=7'b1001111;
        4'h2:a_to_g=7'b0010010;
        4'h3:a_to_g=7'b0000110;
        4'h4:a_to_g=7'b1001100;
        4'h5:a_to_g=7'b0100100;
        4'h6:a_to_g=7'b0100000;
        4'h7:a_to_g=7'b0001111;
        4'h8:a_to_g=7'b0000000;
        4'h9:a_to_g=7'b0000100;
        4'hA:a_to_g=7'b0001000;
        4'hB:a_to_g=7'b1100000;
        4'hC:a_to_g=7'b0110001;
        4'hD:a_to_g=7'b1000010;
        4'hE:a_to_g=7'b0110000;
        4'hF:a_to_g=7'b0111000;
        default:a_to_g=7'b0000001;
    endcase
    always@(*)              //�ı�λ
    begin
        an=4'b1111;
        an[s]=0;
    end
    
    always@(posedge clk)
    begin
        clk_cnt=clk_cnt+1;
    end
endmodule
